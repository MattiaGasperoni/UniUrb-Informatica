//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "it"
//: property prefix = "_GG"
//: property title = "gateCMOS.v"
//: property technology = unit
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] X1;    //: /sn:0 {0}(#:397,371)(397,315){1}
//: {2}(399,313)(433,313)(433,301){3}
//: {4}(397,311)(#:397,259){5}
reg [3:0] C3;    //: /sn:0 {0}(#:1071,371)(1071,305){1}
//: {2}(1073,303)(1102,303)(1102,298){3}
//: {4}(1071,301)(#:1071,253){5}
reg [3:0] C4;    //: /sn:0 {0}(#:1371,256)(1371,306)(1371,306)(1371,316){1}
//: {2}(1373,318)(1408,318)(1408,296){3}
//: {4}(1371,320)(#:1371,376){5}
reg [3:0] X2;    //: /sn:0 {0}(#:688,257)(688,301){1}
//: {2}(690,303)(724,303)(724,295){3}
//: {4}(#:688,305)(688,462)(739,462)(#:739,473){5}
reg [3:0] C2;    //: /sn:0 {0}(#:944,254)(944,309){1}
//: {2}(946,311)(984,311)(984,291){3}
//: {4}(944,313)(#:944,466)(999,466)(#:999,473){5}
reg ENABLE;    //: /sn:0 {0}(89,349)(89,472)(197,472){1}
//: {2}(199,470)(199,352){3}
//: {4}(199,474)(199,515){5}
reg clk;    //: /sn:0 {0}(1331,376)(1331,363)(1297,363){1}
//: {2}(1293,363)(1190,363){3}
//: {4}(1186,363)(1150,363){5}
//: {6}(1146,363)(1032,363){7}
//: {8}(1028,363)(765,363){9}
//: {10}(761,363)(493,363){11}
//: {12}(489,363)(359,363){13}
//: {14}(357,361)(357,371){15}
//: {16}(355,363)(319,363){17}
//: {18}(315,363)(130,363){19}
//: {20}(128,361)(128,352){21}
//: {22}(128,365)(128,515){23}
//: {24}(317,365)(317,713)(700,713){25}
//: {26}(491,365)(491,371){27}
//: {28}(763,365)(763,371){29}
//: {30}(1030,365)(1030,371){31}
//: {32}(1148,365)(1148,441){33}
//: {34}(1150,443)(1189,443)(1189,451){35}
//: {36}(1148,445)(1148,528)(1190,528)(1190,537){37}
//: {38}(1188,365)(1188,371){39}
//: {40}(1295,365)(1295,440){41}
//: {42}(1297,442)(1332,442)(1332,452){43}
//: {44}(1295,444)(1295,527)(1333,527)(1333,537){45}
reg [3:0] X4;    //: /sn:0 {0}(#:1228,371)(1228,308){1}
//: {2}(1230,306)(1266,306)(1266,296){3}
//: {4}(1228,304)(#:1228,256){5}
reg [3:0] C1;    //: /sn:0 {0}(#:531,371)(531,310){1}
//: {2}(533,308)(566,308)(566,297){3}
//: {4}(531,306)(#:531,258){5}
reg [3:0] X3;    //: /sn:0 {0}(#:803,371)(803,304){1}
//: {2}(805,302)(838,302)(838,293){3}
//: {4}(803,300)(#:803,255){5}
wire [7:0] SOMMA;    //: /sn:0 {0}(#:749,733)(749,752){1}
wire [3:0] w58;    //: /sn:0 {0}(#:1072,425)(1072,454)(1039,454)(#:1039,473){1}
wire [3:0] VAL2_2;    //: /sn:0 {0}(#:1021,536)(1021,643)(779,643)(779,674){1}
wire [3:0] VAL1_2;    //: /sn:0 {0}(#:532,424)(532,609)(740,609)(740,674){1}
wire [3:0] w50;    //: /sn:0 {0}(#:804,425)(804,462)(#:779,462)(779,473){1}
wire [3:0] VAL2_1;    //: /sn:0 {0}(#:761,535)(761,674){1}
wire w3;    //: /sn:0 {0}(66,349)(66,596)(167,596){1}
//: {2}(171,596)(331,596){3}
//: {4}(335,596)(697,596){5}
//: {6}(701,596)(959,596)(959,505)(968,505){7}
//: {8}(699,594)(699,504)(708,504){9}
//: {10}(333,598)(333,693)(700,693){11}
//: {12}(169,594)(169,575){13}
wire [3:0] w22;    //: /sn:0 {0}(#:1229,425)(#:1229,451){1}
wire [7:0] TOT;    //: /sn:0 {0}(278,299)(#:278,837)(750,837)(750,822){1}
wire [3:0] MUL4_1;    //: /sn:0 {0}(#:1231,591)(1231,769)(834,769){1}
wire w8;    //: /sn:0 {0}(300,332)(300,788)(668,788){1}
wire [3:0] w11;    //: /sn:0 {0}(#:1372,430)(#:1372,452){1}
wire [3:0] w2;    //: /sn:0 {0}(#:1230,537)(#:1230,505){1}
wire [3:0] VAL1_1;    //: /sn:0 {0}(719,674)(719,628)(#:398,628)(#:398,425){1}
wire [3:0] MUL4_2;    //: /sn:0 {0}(#:1374,591)(1374,806)(834,806){1}
wire [3:0] w5;    //: /sn:0 {0}(#:1373,537)(#:1373,506){1}
//: enddecls

  //: DIP g4 (C2) @(944,244) /sn:0 /w:[ 0 ] /st:10 /dn:1
  //: joint g44 (clk) @(1295, 442) /w:[ 42 41 -1 44 ]
  SReg4 g8 (.clk(clk), .in(C1), .out(VAL1_2));   //: @(477, 372) /sz:(106, 51) /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  //: joint g16 (clk) @(128, 363) /w:[ 19 20 -1 22 ]
  MUX2x4 g47 (.IN0(C2), .IN1(w58), .c(w3), .OUT(VAL2_2));   //: @(969, 474) /sz:(98, 61) /sn:0 /p:[ Ti0>5 Ti1>1 Li0>7 Bo0<0 ]
  //: DIP g3 (C1) @(531,248) /sn:0 /w:[ 5 ] /st:4 /dn:1
  //: joint g17 (w3) @(169, 596) /w:[ 2 12 1 -1 ]
  SReg4 g26 (.in(X4), .clk(clk), .out(w22));   //: @(1174, 372) /sz:(106, 52) /sn:0 /p:[ Ti0>0 Ti1>39 Bo0<0 ]
  //: DIP g2 (X3) @(803,245) /sn:0 /w:[ 5 ] /st:4 /dn:1
  //: joint g23 (C3) @(1071, 303) /w:[ 2 4 -1 1 ]
  //: joint g30 (clk) @(1148, 363) /w:[ 5 -1 6 32 ]
  //: DIP g1 (X2) @(688,247) /sn:0 /w:[ 0 ] /st:5 /dn:1
  //: SWITCH g86 (ENABLE) @(199,339) /sn:0 /R:3 /w:[ 3 ] /st:1 /dn:1
  //: DIP g77 (C4) @(1371,246) /sn:0 /w:[ 0 ] /st:2 /dn:1
  //: joint g24 (clk) @(1030, 363) /w:[ 7 -1 8 30 ]
  SReg4 g29 (.in(w22), .clk(clk), .out(w2));   //: @(1175, 452) /sz:(106, 52) /sn:0 /p:[ Ti0>1 Ti1>35 Bo0<1 ]
  //: LED g60 (X1) @(433,294) /sn:0 /w:[ 3 ] /type:3
  //: joint g51 (clk) @(357, 363) /w:[ 13 14 16 -1 ]
  SReg4 g18 (.in(X3), .clk(clk), .out(w50));   //: @(749, 372) /sz:(106, 52) /sn:0 /p:[ Ti0>0 Ti1>29 Bo0<0 ]
  //: LED g82 (w3) @(66,342) /sn:0 /w:[ 0 ] /type:0
  //: LED g65 (C3) @(1102,291) /sn:0 /w:[ 3 ] /type:3
  MUX2x4 g25 (.IN0(X2), .IN1(w50), .c(w3), .OUT(VAL2_1));   //: @(709, 474) /sz:(98, 60) /sn:0 /p:[ Ti0>5 Ti1>1 Li0>9 Bo0<0 ]
  //: DIP g94 (X4) @(1228,246) /sn:0 /w:[ 5 ] /st:10 /dn:1
  //: joint g10 (C2) @(944, 311) /w:[ 2 1 -1 4 ]
  //: LED g64 (C2) @(984,284) /sn:0 /w:[ 3 ] /type:3
  //: joint g49 (C1) @(531, 308) /w:[ 2 4 -1 1 ]
  SReg4 g6 (.clk(clk), .in(X1), .out(VAL1_1));   //: @(343, 372) /sz:(106, 52) /sn:0 /p:[ Ti0>15 Ti1>0 Bo0<1 ]
  //: joint g50 (clk) @(491, 363) /w:[ 11 -1 12 26 ]
  //: DIP g7 (C3) @(1071,243) /sn:0 /w:[ 5 ] /st:8 /dn:1
  //: joint g9 (X2) @(688, 303) /w:[ 2 1 -1 4 ]
  //: joint g35 (clk) @(1295, 363) /w:[ 1 -1 2 40 ]
  //: joint g31 (C4) @(1371, 318) /w:[ 2 1 -1 4 ]
  SReg4 g22 (.in(C3), .clk(clk), .out(w58));   //: @(1017, 372) /sz:(106, 52) /sn:0 /p:[ Ti0>0 Ti1>31 Bo0<0 ]
  CU g36 (.clk(clk), .enable(ENABLE), .c(w3));   //: @(110, 516) /sz:(122, 58) /sn:0 /p:[ Ti0>23 Ti1>5 Bo0<13 ]
  SReg4 g33 (.in(w11), .clk(clk), .out(w5));   //: @(1318, 453) /sz:(106, 52) /sn:0 /p:[ Ti0>1 Ti1>43 Bo0<1 ]
  //: LED g45 (TOT) @(278,292) /sn:0 /w:[ 0 ] /type:3
  SReg4 g41 (.clk(clk), .in(w2), .out(MUL4_1));   //: @(1176, 538) /sz:(106, 52) /sn:0 /p:[ Ti0>37 Ti1>0 Bo0<0 ]
  //: LED g81 (ENABLE) @(89,342) /sn:0 /w:[ 0 ] /type:0
  //: joint g40 (clk) @(1148, 443) /w:[ 34 33 -1 36 ]
  SReg4 g42 (.clk(clk), .in(w5), .out(MUL4_2));   //: @(1319, 538) /sz:(106, 52) /sn:0 /p:[ Ti0>45 Ti1>0 Bo0<0 ]
  //: LED g12 (w8) @(300,325) /sn:0 /tech:unit /w:[ 0 ] /type:0
  SReg4 g34 (.in(C4), .clk(clk), .out(w11));   //: @(1317, 377) /sz:(106, 52) /sn:0 /p:[ Ti0>5 Ti1>0 Bo0<0 ]
  //: joint g28 (clk) @(1188, 363) /w:[ 3 -1 4 38 ]
  //: joint g46 (X1) @(397, 313) /w:[ 2 4 -1 1 ]
  //: joint g5 (clk) @(317, 363) /w:[ 17 -1 18 24 ]
  //: SWITCH g11 (clk) @(128,339) /sn:0 /R:3 /w:[ 21 ] /st:1 /dn:1
  //: joint g14 (w3) @(333, 596) /w:[ 4 -1 3 10 ]
  MUL_ADD MUL_ADD (.A(VAL1_1), .B(VAL1_2), .C(VAL2_1), .D(VAL2_2), .c(w3), .clk(clk), .S(SOMMA));   //: @(701, 675) /sz:(98, 57) /sn:0 /p:[ Ti0>0 Ti1>1 Ti2>1 Ti3>1 Li0>11 Li1>25 Bo0<0 ]
  //: joint g21 (clk) @(763, 363) /w:[ 9 -1 10 28 ]
  //: LED g61 (C1) @(566,290) /sn:0 /w:[ 3 ] /type:3
  MUL_SUB g19 (.A(SOMMA), .B(MUL4_1), .C(MUL4_2), .Cout(w8), .S(TOT));   //: @(669, 753) /sz:(164, 68) /sn:0 /p:[ Ti0>1 Ri0>1 Ri1>1 Lo0<1 Bo0<1 ]
  //: joint g20 (X3) @(803, 302) /w:[ 2 4 -1 1 ]
  //: LED g78 (X4) @(1266,289) /sn:0 /w:[ 3 ] /type:3
  //: LED g63 (X3) @(838,286) /sn:0 /w:[ 3 ] /type:3
  //: DIP g0 (X1) @(397,249) /sn:0 /w:[ 5 ] /st:10 /dn:1
  //: LED g89 (C4) @(1408,289) /sn:0 /w:[ 3 ] /type:3
  //: joint g27 (X4) @(1228, 306) /w:[ 2 4 -1 1 ]
  //: LED g62 (X2) @(724,288) /sn:0 /w:[ 3 ] /type:3
  //: joint g13 (ENABLE) @(199, 472) /w:[ -1 2 1 4 ]
  //: joint g76 (w3) @(699, 596) /w:[ 6 8 5 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFDls
module FFDls(Y, clk, D);
//: interface  /sz:(40, 40) /bd:[ Li0>D(9/40) Li1>clk(30/40) Ro0<Y(10/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input clk;    //: /sn:0 {0}(189,202)(189,153){1}
//: {2}(191,151)(221,151){3}
//: {4}(189,149)(189,113)(221,113){5}
input D;    //: /sn:0 {0}(157,110)(157,103)(156,103)(156,94){1}
//: {2}(158,92)(221,92){3}
//: {4}(154,92)(139,92){5}
output Y;    //: /sn:0 {0}(470,110)(422,110){1}
wire w3;    //: /sn:0 {0}(437,134)(422,134){1}
wire w0;    //: /sn:0 {0}(301,103)(337,103)(337,109)(347,109){1}
wire w1;    //: /sn:0 {0}(305,162)(337,162)(337,138)(347,138){1}
wire w5;    //: /sn:0 {0}(221,172)(159,172)(159,160){1}
//: enddecls

  //: joint g8 (clk) @(189, 151) /w:[ 2 4 -1 1 ]
  myAND g4 (.in2(w5), .in1(clk), .out(w1));   //: @(222, 141) /sz:(82, 45) /sn:0 /p:[ Li0>0 Li1>3 Ro0<0 ]
  LatchSR g3 (.r(w1), .s(w0), .Y1(w3), .Y(Y));   //: @(348, 101) /sz:(73, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<1 ]
  //: OUT g2 (Y) @(467,110) /sn:0 /w:[ 0 ]
  //: IN g1 (clk) @(189,204) /sn:0 /R:1 /w:[ 0 ]
  myINV g6 (.in(D), .out(w5));   //: @(130, 111) /sz:(52, 48) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  //: joint g7 (D) @(156, 92) /w:[ 2 -1 4 1 ]
  myAND g5 (.in2(clk), .in1(D), .out(w0));   //: @(222, 83) /sz:(78, 44) /sn:0 /p:[ Li0>5 Li1>3 Ro0<0 ]
  //: IN g0 (D) @(137,92) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin myMUX2
module myMUX2(out, c, a, b);
//: interface  /sz:(40, 62) /bd:[ Li0>a(14/62) Li1>b(45/62) Bi0>c(19/40) Ro0<out(29/62) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(166,190)(301,190){1}
output out;    //: /sn:0 {0}(555,131)(523,131){1}
input a;    //: /sn:0 {0}(162,68)(299,68){1}
input c;    //: /sn:0 {0}(301,168)(238,168){1}
//: {2}(236,166)(236,144){3}
//: {4}(236,170)(236,252){5}
wire w7;    //: /sn:0 {0}(392,177)(419,177)(419,144)(434,144){1}
wire w4;    //: /sn:0 {0}(389,76)(418,76)(418,122)(434,122){1}
wire w1;    //: /sn:0 {0}(234,94)(234,89)(299,89){1}
//: enddecls

  //: OUT g8 (out) @(552,131) /sn:0 /w:[ 0 ]
  //: IN g4 (c) @(236,254) /sn:0 /R:1 /w:[ 5 ]
  myNAND g3 (.in1(w4), .in2(w7), .out(out));   //: @(435, 108) /sz:(87, 52) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 ]
  myNAND g2 (.in1(c), .in2(b), .out(w7));   //: @(302, 155) /sz:(89, 50) /sn:0 /p:[ Li0>0 Li1>1 Ro0<0 ]
  myNAND g1 (.in1(a), .in2(w1), .out(w4));   //: @(300, 54) /sz:(88, 51) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: IN g6 (a) @(160,68) /sn:0 /w:[ 0 ]
  //: IN g7 (b) @(164,190) /sn:0 /w:[ 0 ]
  //: joint g5 (c) @(236, 168) /w:[ 1 2 -1 4 ]
  myINV g0 (.in(c), .out(w1));   //: @(215, 95) /sz:(45, 48) /R:1 /sn:0 /p:[ Bi0>3 To0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin CU
module CU(clk, enable, c);
//: interface  /sz:(112, 58) /bd:[ Ti0>enable(79/112) Ti1>clk(8/112) Bo0<c(20/112) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input enable;    //: /sn:0 {0}(180,164)(244,164){1}
input clk;    //: /sn:0 {0}(388,196)(370,196)(370,269)(348,269){1}
output c;    //: /sn:0 {0}(502,190)(502,173){1}
//: {2}(504,171)(458,171)(458,171)(579,171){3}
//: {4}(500,171)(454,171){5}
wire w4;    //: /sn:0 {0}(505,232)(505,239)(230,239)(230,184)(244,184){1}
wire w1;    //: /sn:0 {0}(321,170)(388,170){1}
//: enddecls

  myINV g4 (.in(c), .out(w4));   //: @(477, 191) /sz:(49, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  //: IN g3 (clk) @(346,269) /sn:0 /w:[ 1 ]
  //: joint g6 (c) @(502, 171) /w:[ 2 -1 4 1 ]
  myAND g9 (.in2(w4), .in1(enable), .out(w1));   //: @(245, 155) /sz:(75, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: IN g7 (enable) @(178,164) /sn:0 /w:[ 0 ]
  //: OUT g5 (c) @(576,171) /sn:0 /w:[ 3 ]
  FFDet g0 (.D(w1), .clk(clk), .Y(c));   //: @(389, 161) /sz:(64, 47) /sn:0 /p:[ Li0>1 Li1>0 Ro0<5 ]

endmodule
//: /netlistEnd

//: /netlistBegin RCA8
module RCA8(A, Cout, Cin, B, S);
//: interface  /sz:(125, 44) /bd:[ Ti0>A[7:0](29/125) Ti1>B[7:0](93/125) Ri0>Cin(21/44) Lo0<Cout(23/44) Bo0<S[7:0](60/125) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:-300,51)(-208,51){1}
//: {2}(-207,51)(-105,51){3}
//: {4}(-104,51)(-9,51){5}
//: {6}(-8,51)(84,51){7}
//: {8}(85,51)(175,51){9}
//: {10}(176,51)(266,51){11}
//: {12}(267,51)(359,51){13}
//: {14}(360,51)(455,51){15}
//: {16}(456,51)(501,51){17}
input [7:0] A;    //: /sn:0 {0}(#:-300,29)(-242,29){1}
//: {2}(-241,29)(-139,29){3}
//: {4}(-138,29)(-43,29){5}
//: {6}(-42,29)(51,29){7}
//: {8}(52,29)(143,29){9}
//: {10}(144,29)(233,29){11}
//: {12}(234,29)(325,29){13}
//: {14}(326,29)(423,29){15}
//: {16}(424,29)(491,29){17}
input Cin;    //: /sn:0 {0}(501,113)(478,113){1}
output Cout;    //: /sn:0 {0}(-283,105)(-261,105){1}
output [7:0] S;    //: /sn:0 {0}(#:103,209)(103,273){1}
wire w16;    //: /sn:0 {0}(33,108)(15,108){1}
wire w13;    //: /sn:0 {0}(108,203)(108,182)(160,182)(160,140){1}
wire w6;    //: /sn:0 {0}(456,55)(456,86){1}
wire w7;    //: /sn:0 {0}(383,112)(406,112){1}
wire w34;    //: /sn:0 {0}(-241,33)(-241,79){1}
wire w25;    //: /sn:0 {0}(360,55)(360,85){1}
wire w4;    //: /sn:0 {0}(118,203)(118,186)(250,186)(250,141){1}
wire w22;    //: /sn:0 {0}(-158,106)(-184,106){1}
wire w3;    //: /sn:0 {0}(215,110)(198,110){1}
wire w0;    //: /sn:0 {0}(234,33)(234,85){1}
wire w20;    //: /sn:0 {0}(-104,55)(-104,80){1}
wire w30;    //: /sn:0 {0}(85,55)(85,83){1}
wire w29;    //: /sn:0 {0}(52,33)(52,83){1}
wire w19;    //: /sn:0 {0}(-138,33)(-138,80){1}
wire w18;    //: /sn:0 {0}(88,203)(88,185)(-26,185)(-26,140){1}
wire w12;    //: /sn:0 {0}(126,109)(107,109){1}
wire w23;    //: /sn:0 {0}(-122,140)(-122,189)(78,189)(78,203){1}
wire w10;    //: /sn:0 {0}(176,55)(176,84){1}
wire w24;    //: /sn:0 {0}(326,33)(326,85){1}
wire w1;    //: /sn:0 {0}(267,55)(267,85){1}
wire w8;    //: /sn:0 {0}(138,203)(138,193)(440,193)(440,145){1}
wire w17;    //: /sn:0 {0}(-61,107)(-81,107){1}
wire w33;    //: /sn:0 {0}(98,203)(98,182)(68,182)(68,141){1}
wire w35;    //: /sn:0 {0}(-207,55)(-207,79){1}
wire w28;    //: /sn:0 {0}(342,144)(342,190)(128,190)(128,203){1}
wire w14;    //: /sn:0 {0}(-42,33)(-42,81){1}
wire w2;    //: /sn:0 {0}(307,111)(289,111){1}
wire w15;    //: /sn:0 {0}(-8,55)(-8,81){1}
wire w5;    //: /sn:0 {0}(424,33)(424,86){1}
wire w38;    //: /sn:0 {0}(-225,139)(-225,192)(68,192)(68,203){1}
wire w9;    //: /sn:0 {0}(144,33)(144,84){1}
//: enddecls

  FA g4 (.B(w20), .A(w19), .Cin(w17), .Cout(w22), .S(w23));   //: @(-157, 81) /sz:(75, 58) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: IN g8 (A) @(-302,29) /sn:0 /w:[ 0 ]
  FA g3 (.B(w15), .A(w14), .Cin(w16), .Cout(w17), .S(w18));   //: @(-60, 82) /sz:(74, 57) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  assign w24 = A[1]; //: TAP g16 @(326,27) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  assign w19 = A[6]; //: TAP g17 @(-138,27) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: OUT g26 (Cout) @(-280,105) /sn:0 /R:2 /w:[ 0 ]
  FA g2 (.B(w10), .A(w9), .Cin(w3), .Cout(w12), .S(w13));   //: @(127, 85) /sz:(70, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: IN g30 (Cin) @(503,113) /sn:0 /R:2 /w:[ 0 ]
  assign w34 = A[7]; //: TAP g23 @(-241,27) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w35 = B[7]; //: TAP g24 @(-207,49) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  FA g1 (.B(w6), .A(w5), .Cin(Cin), .Cout(w7), .S(w8));   //: @(407, 87) /sz:(70, 57) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  assign w20 = B[6]; //: TAP g18 @(-104,49) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign w5 = A[0]; //: TAP g10 @(424,27) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  assign w25 = B[1]; //: TAP g25 @(360,49) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  FA g6 (.B(w30), .A(w29), .Cin(w12), .Cout(w16), .S(w33));   //: @(34, 84) /sz:(72, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  FA g7 (.B(w35), .A(w34), .Cin(w22), .Cout(Cout), .S(w38));   //: @(-260, 80) /sz:(75, 58) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  //: IN g9 (B) @(-302,51) /sn:0 /w:[ 0 ]
  assign w1 = B[2]; //: TAP g22 @(267,49) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  assign w29 = A[4]; //: TAP g12 @(52,27) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign S = {w38, w23, w18, w33, w13, w4, w28, w8}; //: CONCAT g28  @(103,208) /sn:0 /R:3 /w:[ 0 1 1 0 0 0 0 1 0 ] /dr:1 /tp:0 /drp:1
  FA g5 (.B(w25), .A(w24), .Cin(w7), .Cout(w2), .S(w28));   //: @(308, 86) /sz:(74, 57) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  assign w6 = B[0]; //: TAP g11 @(456,49) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  assign w9 = A[3]; //: TAP g14 @(144,27) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  assign w15 = B[5]; //: TAP g19 @(-8,49) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w10 = B[3]; //: TAP g21 @(176,49) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  assign w30 = B[4]; //: TAP g20 @(85,49) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  FA g0 (.B(w1), .A(w0), .Cin(w2), .Cout(w3), .S(w4));   //: @(216, 86) /sz:(72, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  assign w14 = A[5]; //: TAP g15 @(-42,27) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: OUT g27 (S) @(103,270) /sn:0 /R:3 /w:[ 1 ]
  assign w0 = A[2]; //: TAP g13 @(234,27) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin SUB8
module SUB8(Cin, B, A, S, Cout);
//: interface  /sz:(96, 40) /bd:[ Ti0>B[7:0](51/96) Ti1>A[7:0](21/96) Ri0>Cin(22/40) Lo0<Cout(22/40) Bo0<S[7:0](43/96) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:353,-13)(353,47){1}
input [7:0] A;    //: /sn:0 {0}(#:290,-13)(#:290,147){1}
input Cin;    //: /sn:0 {0}(442,54)(442,169)(387,169){1}
output Cout;    //: /sn:0 {0}(149,66)(149,103){1}
output [7:0] S;    //: /sn:0 {0}(#:321,248)(#:321,193){1}
wire w0;    //: /sn:0 {0}(260,171)(150,171)(150,155){1}
wire [7:0] w1;    //: /sn:0 {0}(354,99)(#:354,147){1}
//: enddecls

  //: IN g4 (Cin) @(442,52) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  //: IN g3 (B) @(353,-15) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  //: IN g2 (A) @(290,-15) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  RCA8 g1 (.A(A), .B(w1), .Cin(Cin), .Cout(w0), .S(S));   //: @(261, 148) /sz:(125, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: OUT g6 (S) @(321,245) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  myINV g7 (.in(w0), .out(Cout));   //: @(125, 104) /sz:(49, 50) /R:1 /sn:0 /p:[ Bi0>1 To0<1 ]
  //: OUT g5 (Cout) @(149,69) /sn:0 /R:1 /tech:unit /w:[ 0 ]
  myINV8 g0 (.IN(B), .OUT(w1));   //: @(327, 48) /sz:(53, 50) /sn:0 /p:[ Ti0>1 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myINV8
module myINV8(IN, OUT);
//: interface  /sz:(53, 50) /bd:[ Ti0>IN[7:0](25/53) Bo0<OUT[7:0](27/53) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output [7:0] OUT;    //: /sn:0 {0}(#:591,86)(627,86){1}
input [7:0] IN;    //: /sn:0 {0}(#:174,-70)(197,-70)(197,-47){1}
//: {2}(197,-46)(197,2){3}
//: {4}(197,3)(197,51){5}
//: {6}(197,52)(197,101){7}
//: {8}(197,102)(197,149){9}
//: {10}(197,150)(197,199){11}
//: {12}(197,200)(197,249){13}
//: {14}(197,250)(197,299){15}
//: {16}(197,300)(197,323){17}
wire w13;    //: /sn:0 {0}(585,101)(518,101)(518,198)(371,198){1}
wire w6;    //: /sn:0 {0}(287,52)(201,52){1}
wire w7;    //: /sn:0 {0}(370,50)(500,50)(500,71)(585,71){1}
wire w4;    //: /sn:0 {0}(287,102)(201,102){1}
wire w0;    //: /sn:0 {0}(287,-47)(209,-47)(209,-46)(201,-46){1}
wire w3;    //: /sn:0 {0}(370,1)(510,1)(510,61)(585,61){1}
wire w12;    //: /sn:0 {0}(287,200)(201,200){1}
wire w10;    //: /sn:0 {0}(287,300)(201,300){1}
wire w1;    //: /sn:0 {0}(369,-49)(554,-49)(554,51)(585,51){1}
wire w8;    //: /sn:0 {0}(287,250)(201,250){1}
wire w14;    //: /sn:0 {0}(287,150)(201,150){1}
wire w11;    //: /sn:0 {0}(373,298)(547,298)(547,121)(585,121){1}
wire w2;    //: /sn:0 {0}(287,3)(201,3){1}
wire w15;    //: /sn:0 {0}(370,148)(511,148)(511,91)(585,91){1}
wire w5;    //: /sn:0 {0}(585,81)(500,81)(500,100)(370,100){1}
wire w9;    //: /sn:0 {0}(585,111)(528,111)(528,248)(372,248){1}
//: enddecls

  myINV g8 (.in(w14), .out(w15));   //: @(288, 131) /sz:(81, 42) /sn:0 /p:[ Li0>0 Ro0<0 ]
  myINV g4 (.in(w6), .out(w7));   //: @(288, 33) /sz:(81, 42) /sn:0 /p:[ Li0>0 Ro0<0 ]
  assign w12 = IN[5]; //: TAP g16 @(195,200) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  myINV g3 (.in(w4), .out(w5));   //: @(288, 83) /sz:(81, 42) /sn:0 /p:[ Li0>0 Ro0<1 ]
  assign w8 = IN[6]; //: TAP g17 @(195,250) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  myINV g2 (.in(w2), .out(w3));   //: @(288, -17) /sz:(81, 43) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: IN g1 (IN) @(172,-70) /sn:0 /w:[ 0 ]
  assign w10 = IN[7]; //: TAP g18 @(195,300) /sn:0 /R:2 /w:[ 1 16 15 ] /ss:1
  assign OUT = {w11, w9, w13, w15, w5, w7, w3, w1}; //: CONCAT g10  @(590,86) /sn:0 /w:[ 0 1 0 0 1 0 1 1 1 ] /dr:1 /tp:0 /drp:1
  myINV g6 (.in(w10), .out(w11));   //: @(288, 281) /sz:(84, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: OUT g9 (OUT) @(624,86) /sn:0 /w:[ 1 ]
  myINV g7 (.in(w12), .out(w13));   //: @(288, 181) /sz:(82, 40) /sn:0 /p:[ Li0>0 Ro0<1 ]
  assign w2 = IN[1]; //: TAP g12 @(195,3) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  assign w4 = IN[3]; //: TAP g14 @(195,102) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  assign w0 = IN[0]; //: TAP g11 @(195,-46) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  myINV g5 (.in(w8), .out(w9));   //: @(288, 231) /sz:(83, 40) /sn:0 /p:[ Li0>0 Ro0<1 ]
  assign w14 = IN[4]; //: TAP g15 @(195,150) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  myINV g0 (.in(w0), .out(w1));   //: @(288, -67) /sz:(80, 44) /sn:0 /p:[ Li0>0 Ro0<0 ]
  assign w6 = IN[2]; //: TAP g13 @(195,52) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin LatchSR
module LatchSR(Y1, Y, r, s);
//: interface  /sz:(40, 40) /bd:[ Li0>s(7/40) Li1>r(31/40) Ro0<Y(8/40) Ro1<Y1(28/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input r;    //: /sn:0 {0}(133,158)(224,158){1}
input s;    //: /sn:0 {0}(132,61)(223,61){1}
output Y1;    //: /sn:0 {0}(224,135)(198,135)(198,114)(341,114)(341,75){1}
//: {2}(343,73)(383,73)(383,76)(410,76){3}
//: {4}(339,73)(313,73){5}
output Y;    //: /sn:0 {0}(315,149)(344,149){1}
//: {2}(348,149)(376,149)(376,148)(415,148){3}
//: {4}(346,147)(346,106)(198,106)(198,82)(223,82){5}
//: enddecls

  myNOR g4 (.in2(Y), .in1(s), .out(Y1));   //: @(224, 50) /sz:(88, 50) /sn:0 /p:[ Li0>5 Li1>1 Ro0<5 ]
  //: OUT g3 (Y1) @(407,76) /sn:0 /w:[ 3 ]
  //: OUT g2 (Y) @(412,148) /sn:0 /w:[ 3 ]
  //: IN g1 (r) @(131,158) /sn:0 /w:[ 0 ]
  //: joint g6 (Y) @(346, 149) /w:[ 2 4 1 -1 ]
  //: joint g7 (Y1) @(341, 73) /w:[ 2 -1 4 1 ]
  myNOR g5 (.in2(r), .in1(Y1), .out(Y));   //: @(225, 124) /sz:(89, 53) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  //: IN g0 (s) @(130,61) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myNAND
module myNAND(out, in2, in1);
//: interface  /sz:(40, 40) /bd:[ Li0>in2(28/40) Li1>in1(11/40) Ro0<out(18/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
supply1 w0;    //: /sn:0 {0}(250,34)(250,42)(251,42)(251,52){1}
//: {2}(253,54)(304,54)(304,88){3}
//: {4}(249,54)(215,54)(215,73){5}
input in1;    //: /sn:0 {0}(121,82)(167,82){1}
//: {2}(171,82)(188,82)(188,81)(201,81){3}
//: {4}(169,84)(169,178)(241,178){5}
supply0 w1;    //: /sn:0 {0}(255,238)(255,278){1}
output out;    //: /sn:0 {0}(255,170)(255,148){1}
//: {2}(257,146)(405,146){3}
//: {4}(255,144)(255,123){5}
//: {6}(257,121)(304,121)(304,105){7}
//: {8}(253,121)(215,121)(215,90){9}
input in2;    //: /sn:0 {0}(121,96)(154,96){1}
//: {2}(158,96)(290,96){3}
//: {4}(156,98)(156,229)(241,229){5}
wire w9;    //: /sn:0 {0}(255,187)(255,221){1}
//: enddecls

  //: GROUND g4 (w1) @(255,284) /sn:0 /w:[ 1 ]
  _GGNMOS #(2, 1) g8 (.Z(w9), .S(w1), .G(in2));   //: @(249,229) /sn:0 /w:[ 1 0 5 ]
  //: VDD g3 (w0) @(261,34) /sn:0 /w:[ 0 ]
  //: OUT g2 (out) @(402,146) /sn:0 /w:[ 3 ]
  //: IN g1 (in2) @(119,96) /sn:0 /w:[ 0 ]
  //: joint g10 (w0) @(251, 54) /w:[ 2 1 4 -1 ]
  _GGPMOS #(2, 1) g6 (.Z(out), .S(w0), .G(in2));   //: @(298,96) /sn:0 /w:[ 7 3 3 ]
  _GGNMOS #(2, 1) g7 (.Z(out), .S(w9), .G(in1));   //: @(249,178) /sn:0 /w:[ 0 0 5 ]
  //: joint g9 (out) @(255, 121) /w:[ 6 -1 8 5 ]
  //: joint g12 (in2) @(156, 96) /w:[ 2 -1 1 4 ]
  _GGPMOS #(2, 1) g5 (.Z(out), .S(w0), .G(in1));   //: @(209,81) /sn:0 /w:[ 9 5 3 ]
  //: joint g11 (in1) @(169, 82) /w:[ 2 -1 1 4 ]
  //: IN g0 (in1) @(119,82) /sn:0 /w:[ 0 ]
  //: joint g13 (out) @(255, 146) /w:[ 2 4 -1 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin HA
module HA(Cout, B, S, A);
//: interface  /sz:(57, 57) /bd:[ Ti0>B(39/57) Ti1>A(12/57) Lo0<Cout(28/57) Bo0<S(28/57) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(77,149)(89,149)(89,148)(136,148){1}
//: {2}(138,146)(138,104)(226,104)(226,89)(277,89){3}
//: {4}(138,150)(138,152)(148,152){5}
input A;    //: /sn:0 {0}(86,75)(112,75){1}
//: {2}(116,75)(140,75){3}
//: {4}(114,77)(114,111)(228,111)(228,124)(264,124)(264,135)(278,135){5}
output Cout;    //: /sn:0 {0}(369,209)(544,209){1}
output S;    //: /sn:0 {0}(509,118)(552,118){1}
wire w6;    //: /sn:0 {0}(367,76)(406,76)(406,110)(416,110){1}
wire w3;    //: /sn:0 {0}(278,197)(255,197)(255,152){1}
//: {2}(257,150)(265,150)(265,155)(278,155){3}
//: {4}(253,150)(230,150){5}
wire w1;    //: /sn:0 {0}(278,217)(236,217)(236,76){1}
//: {2}(238,74)(264,74)(264,67)(277,67){3}
//: {4}(234,74)(221,74){5}
wire w9;    //: /sn:0 {0}(366,144)(406,144)(406,130)(416,130){1}
//: enddecls

  myNAND g4 (.in2(w9), .in1(w6), .out(S));   //: @(417, 97) /sz:(91, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: OUT g8 (Cout) @(541,209) /sn:0 /w:[ 1 ]
  myNAND g3 (.in2(w3), .in1(A), .out(w9));   //: @(279, 123) /sz:(86, 47) /sn:0 /p:[ Li0>3 Li1>5 Ro0<0 ]
  myNAND g2 (.in2(B), .in1(w1), .out(w6));   //: @(278, 54) /sz:(88, 50) /sn:0 /p:[ Li0>3 Li1>3 Ro0<0 ]
  myINV g1 (.in(B), .out(w3));   //: @(149, 131) /sz:(80, 45) /sn:0 /p:[ Li0>5 Ro0<5 ]
  //: joint g10 (B) @(138, 148) /w:[ -1 2 1 4 ]
  //: IN g6 (B) @(75,149) /sn:0 /w:[ 0 ]
  //: OUT g7 (S) @(549,118) /sn:0 /w:[ 1 ]
  //: joint g9 (A) @(114, 75) /w:[ 2 -1 1 4 ]
  //: joint g12 (w3) @(255, 150) /w:[ 2 -1 4 1 ]
  //: IN g5 (A) @(84,75) /sn:0 /w:[ 0 ]
  myNOR g11 (.in1(w3), .in2(w1), .out(Cout));   //: @(279, 187) /sz:(89, 47) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  myINV g0 (.in(A), .out(w1));   //: @(141, 57) /sz:(79, 41) /sn:0 /p:[ Li0>3 Ro0<5 ]
  //: joint g13 (w1) @(236, 74) /w:[ 2 -1 4 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin myEXOR
module myEXOR(out, B, A);
//: interface  /sz:(40, 40) /bd:[ Li0>B(26/40) Li1>A(8/40) Ro0<out(20/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(235,98)(206,98)(206,117)(106,117)(106,151){1}
//: {2}(104,153)(68,153){3}
//: {4}(106,155)(106,180)(112,180){5}
input A;    //: /sn:0 {0}(235,147)(203,147)(203,130)(94,130)(94,66){1}
//: {2}(96,64)(113,64){3}
//: {4}(92,64)(68,64){5}
output out;    //: /sn:0 {0}(456,120)(488,120){1}
wire w6;    //: /sn:0 {0}(329,85)(357,85)(357,113)(365,113){1}
wire w3;    //: /sn:0 {0}(204,179)(224,179)(224,171)(235,171){1}
wire w1;    //: /sn:0 {0}(204,61)(225,61)(225,76)(235,76){1}
wire w9;    //: /sn:0 {0}(331,156)(357,156)(357,131)(365,131){1}
//: enddecls

  myINV g4 (.in(B), .out(w3));   //: @(113, 158) /sz:(90, 48) /sn:0 /p:[ Li0>5 Ro0<0 ]
  //: joint g8 (A) @(94, 64) /w:[ 2 -1 4 1 ]
  myINV g3 (.in(A), .out(w1));   //: @(114, 39) /sz:(89, 53) /sn:0 /p:[ Li0>3 Ro0<0 ]
  //: OUT g2 (out) @(485,120) /sn:0 /w:[ 1 ]
  //: IN g1 (B) @(66,153) /sn:0 /w:[ 3 ]
  myNAND g6 (.in2(w3), .in1(A), .out(w9));   //: @(236, 132) /sz:(94, 56) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  myNAND g7 (.in2(w9), .in1(w6), .out(out));   //: @(366, 101) /sz:(89, 44) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: joint g9 (B) @(106, 153) /w:[ -1 1 2 4 ]
  myNAND g5 (.in2(B), .in1(w1), .out(w6));   //: @(236, 62) /sz:(92, 52) /sn:0 /p:[ Li0>0 Li1>1 Ro0<0 ]
  //: IN g0 (A) @(66,64) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFDet
module FFDet(Y, clk, D);
//: interface  /sz:(40, 40) /bd:[ Li0>D(8/40) Li1>clk(30/40) Ro0<Y(9/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input clk;    //: /sn:0 {0}(231,143)(244,143){1}
//: {2}(246,141)(246,97)(257,97){3}
//: {4}(246,145)(246,189){5}
input D;    //: /sn:0 {0}(93,75)(160,75){1}
output Y;    //: /sn:0 {0}(320,77)(364,77){1}
wire w1;    //: /sn:0 {0}(147,139)(132,139)(132,96)(160,96){1}
wire w2;    //: /sn:0 {0}(220,76)(257,76){1}
//: enddecls

  FFDls g4 (.clk(clk), .D(w2), .Y(Y));   //: @(258, 67) /sz:(61, 40) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 ]
  FFDls g3 (.clk(w1), .D(D), .Y(w2));   //: @(161, 66) /sz:(58, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: OUT g2 (Y) @(361,77) /sn:0 /w:[ 1 ]
  //: IN g1 (clk) @(246,191) /sn:0 /R:1 /w:[ 5 ]
  //: joint g6 (clk) @(246, 143) /w:[ -1 2 1 4 ]
  myINV g5 (.in(clk), .out(w1));   //: @(148, 117) /sz:(82, 52) /R:2 /sn:0 /p:[ Ri0>0 Lo0<0 ]
  //: IN g0 (D) @(91,75) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myNOR
module myNOR(out, in2, in1);
//: interface  /sz:(40, 40) /bd:[ Li0>in1(9/40) Li1>in2(26/40) Ro0<out(19/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
supply1 w0;    //: /sn:0 {0}(257,42)(257,78){1}
input in1;    //: /sn:0 {0}(144,126)(202,126){1}
//: {2}(204,124)(204,86)(243,86){3}
//: {4}(204,128)(204,203)(283,203){5}
supply0 w1;    //: /sn:0 {0}(253,263)(253,238){1}
//: {2}(255,236)(297,236)(297,212){3}
//: {4}(251,236)(230,236)(230,222){5}
output out;    //: /sn:0 {0}(256,149)(256,160){1}
//: {2}(258,162)(268,162)(268,150)(403,150){3}
//: {4}(256,164)(256,178){5}
//: {6}(258,180)(297,180)(297,195){7}
//: {8}(254,180)(230,180)(230,205){9}
input in2;    //: /sn:0 {0}(140,172)(188,172){1}
//: {2}(190,170)(190,140)(242,140){3}
//: {4}(190,174)(190,213)(216,213){5}
wire w2;    //: /sn:0 {0}(256,132)(256,117)(257,117)(257,95){1}
//: enddecls

  _GGNMOS #(2, 1) g8 (.Z(out), .S(w1), .G(in1));   //: @(291,203) /sn:0 /w:[ 7 3 5 ]
  //: GROUND g4 (w1) @(253,269) /sn:0 /w:[ 0 ]
  //: VDD g3 (w0) @(268,42) /sn:0 /w:[ 0 ]
  //: OUT g2 (out) @(400,150) /sn:0 /w:[ 3 ]
  //: IN g1 (in2) @(138,172) /sn:0 /w:[ 0 ]
  //: joint g10 (w1) @(253, 236) /w:[ 2 -1 4 1 ]
  _GGPMOS #(2, 1) g6 (.Z(out), .S(w2), .G(in2));   //: @(250,140) /sn:0 /w:[ 0 0 3 ]
  //: joint g9 (out) @(256, 180) /w:[ 6 5 8 -1 ]
  _GGNMOS #(2, 1) g7 (.Z(out), .S(w1), .G(in2));   //: @(224,213) /sn:0 /w:[ 9 5 5 ]
  //: joint g12 (in2) @(190, 172) /w:[ -1 2 1 4 ]
  //: joint g11 (in1) @(204, 126) /w:[ -1 2 1 4 ]
  _GGPMOS #(2, 1) g5 (.Z(w2), .S(w0), .G(in1));   //: @(251,86) /sn:0 /w:[ 1 1 3 ]
  //: IN g0 (in1) @(142,126) /sn:0 /w:[ 0 ]
  //: joint g13 (out) @(256, 162) /w:[ 2 1 -1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin RCA4
module RCA4(A, Cout, Cin, B, S);
//: interface  /sz:(98, 40) /bd:[ Ti0>B[3:0](70/98) Ti1>A[3:0](28/98) Ri0>Cin(20/40) Lo0<Cout(21/40) Bo0<S[7:0](50/98) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] B;    //: /sn:0 {0}(#:-92,42)(84,42){1}
//: {2}(85,42)(176,42){3}
//: {4}(177,42)(262,42){5}
//: {6}(263,42)(352,42){7}
//: {8}(353,42)(375,42){9}
input [3:0] A;    //: /sn:0 {0}(#:-91,20)(58,20){1}
//: {2}(59,20)(150,20){3}
//: {4}(151,20)(236,20){5}
//: {6}(237,20)(325,20){7}
//: {8}(326,20)(372,20){9}
input Cin;    //: /sn:0 {0}(527,92)(395,92)(395,95)(369,95){1}
output Cout;    //: /sn:0 {0}(-82,97)(45,97){1}
output [7:0] S;    //: /sn:0 {0}(#:151,210)(151,242)(150,242)(150,274){1}
wire w13;    //: /sn:0 {0}(136,204)(136,178)(72,178)(72,128){1}
wire w6;    //: /sn:0 {0}(353,46)(353,54)(352,54)(352,69){1}
wire w7;    //: /sn:0 {0}(278,97)(291,97)(291,94)(312,94){1}
wire w25;    //: /sn:0 {0}(263,46)(263,55)(261,55)(261,71){1}
wire w4;    //: /sn:0 {0}(146,204)(146,181)(163,181)(163,126){1}
wire w3;    //: /sn:0 {0}(136,95)(103,95)(103,98)(102,98){1}
wire w0;    //: /sn:0 {0}(151,24)(151,70){1}
wire w10;    //: /sn:0 {0}(85,46)(85,72){1}
wire w24;    //: /sn:0 {0}(237,24)(237,48)(236,48)(236,71){1}
wire w1;    //: /sn:0 {0}(177,46)(177,54)(176,54)(176,70){1}
wire w8;    //: /sn:0 {0}(166,204)(166,194)(339,194)(339,125){1}
wire w28;    //: /sn:0 {0}(248,127)(248,186)(156,186)(156,204){1}
wire w2;    //: /sn:0 {0}(221,96)(193,96){1}
wire w5;    //: /sn:0 {0}(326,24)(326,54)(327,54)(327,69){1}
wire w9;    //: /sn:0 {0}(59,24)(59,32)(60,32)(60,72){1}
//: enddecls

  //: IN g8 (A) @(-93,20) /sn:0 /w:[ 0 ]
  assign w24 = A[1]; //: TAP g16 @(237,18) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: OUT g26 (Cout) @(-79,97) /sn:0 /R:2 /w:[ 0 ]
  FA g2 (.B(w10), .A(w9), .Cin(w3), .Cout(Cout), .S(w13));   //: @(46, 73) /sz:(55, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  //: IN g30 (Cin) @(529,92) /sn:0 /R:2 /w:[ 0 ]
  FA g1 (.B(w6), .A(w5), .Cin(Cin), .Cout(w7), .S(w8));   //: @(313, 70) /sz:(55, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  assign w5 = A[0]; //: TAP g10 @(326,18) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w25 = B[1]; //: TAP g25 @(263,40) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: IN g9 (B) @(-94,42) /sn:0 /w:[ 0 ]
  assign w1 = B[2]; //: TAP g22 @(177,40) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign S = {w13, w4, w28, w8}; //: CONCAT g28  @(151,209) /sn:0 /R:3 /w:[ 0 0 0 1 0 ] /dr:1 /tp:0 /drp:1
  FA g5 (.B(w25), .A(w24), .Cin(w7), .Cout(w2), .S(w28));   //: @(222, 72) /sz:(55, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  assign w6 = B[0]; //: TAP g11 @(353,40) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w9 = A[3]; //: TAP g14 @(59,18) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w10 = B[3]; //: TAP g21 @(85,40) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  FA g0 (.B(w1), .A(w0), .Cin(w2), .Cout(w3), .S(w4));   //: @(137, 71) /sz:(55, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: OUT g27 (S) @(150,271) /sn:0 /R:3 /w:[ 1 ]
  assign w0 = A[2]; //: TAP g13 @(151,18) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin myAND
module myAND(out, in2, in1);
//: interface  /sz:(40, 40) /bd:[ Li0>in1(9/40) Li1>in2(28/40) Ro0<out(19/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(229,142)(159,142){1}
output out;    //: /sn:0 {0}(463,152)(536,152){1}
input in2;    //: /sn:0 {0}(153,171)(205,171)(205,171)(229,171){1}
wire w2;    //: /sn:0 {0}(378,154)(321,154){1}
//: enddecls

  myINV g4 (.in(w2), .out(out));   //: @(379, 130) /sz:(83, 51) /sn:0 /p:[ Li0>0 Ro0<0 ]
  myNAND g3 (.in1(in1), .in2(in2), .out(w2));   //: @(230, 124) /sz:(90, 68) /sn:0 /p:[ Li0>0 Li1>1 Ro0<1 ]
  //: OUT g2 (out) @(533,152) /sn:0 /w:[ 1 ]
  //: IN g1 (in2) @(151,171) /sn:0 /w:[ 0 ]
  //: IN g0 (in1) @(157,142) /sn:0 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin myINV
module myINV(in, out);
//: interface  /sz:(40, 40) /bd:[ Li0>in(19/40) Ro0<out(17/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
supply1 w6;    //: /sn:0 {0}(281,81)(281,115){1}
supply0 w7;    //: /sn:0 {0}(281,190)(281,233){1}
input in;    //: /sn:0 {0}(179,150)(250,150){1}
//: {2}(252,148)(252,123)(267,123){3}
//: {4}(252,152)(252,181)(267,181){5}
output out;    //: /sn:0 {0}(281,132)(281,145){1}
//: {2}(283,147)(330,147)(330,121)(364,121){3}
//: {4}(281,149)(281,173){5}
//: enddecls

  //: IN g4 (in) @(177,150) /sn:0 /w:[ 0 ]
  //: GROUND g3 (w7) @(281,239) /sn:0 /w:[ 1 ]
  //: VDD g2 (w6) @(292,81) /sn:0 /w:[ 0 ]
  _GGNMOS #(2, 1) g1 (.Z(out), .S(w7), .G(in));   //: @(275,181) /sn:0 /w:[ 5 0 5 ]
  //: OUT g6 (out) @(361,121) /sn:0 /w:[ 3 ]
  //: joint g7 (out) @(281, 147) /w:[ 2 1 -1 4 ]
  //: joint g5 (in) @(252, 150) /w:[ -1 2 1 4 ]
  _GGPMOS #(2, 1) g0 (.Z(out), .S(w6), .G(in));   //: @(275,123) /sn:0 /w:[ 0 1 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin SReg8
module SReg8(out, clk, in);
//: interface  /sz:(88, 48) /bd:[ Ti0>in[7:0](41/88) Ti1>clk(10/88) Bo0<out[7:0](42/88) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] in;    //: /sn:0 {0}(#:160,39)(160,77){1}
//: {2}(160,78)(160,124){3}
//: {4}(160,125)(160,172){5}
//: {6}(160,173)(160,222){7}
//: {8}(160,223)(160,277){9}
//: {10}(160,278)(160,330){11}
//: {12}(160,331)(160,385){13}
//: {14}(160,386)(160,440){15}
//: {16}(160,441)(160,500){17}
input clk;    //: /sn:0 {0}(251,102)(208,102)(208,147){1}
//: {2}(210,149)(251,149){3}
//: {4}(208,151)(208,194){5}
//: {6}(210,196)(251,196){7}
//: {8}(208,198)(208,246){9}
//: {10}(210,248)(252,248){11}
//: {12}(208,250)(208,298){13}
//: {14}(210,300)(252,300){15}
//: {16}(208,302)(208,353){17}
//: {18}(210,355)(252,355){19}
//: {20}(208,357)(208,408){21}
//: {22}(210,410)(251,410){23}
//: {24}(208,412)(208,463){25}
//: {26}(210,465)(251,465){27}
//: {28}(208,467)(208,510){29}
output [7:0] out;    //: /sn:0 {0}(#:812,256)(#:741,256){1}
wire w16;    //: /sn:0 {0}(318,224)(686,224)(686,251)(735,251){1}
wire w6;    //: /sn:0 {0}(318,387)(708,387)(708,281)(735,281){1}
wire w13;    //: /sn:0 {0}(164,441)(251,441){1}
wire w7;    //: /sn:0 {0}(252,331)(164,331){1}
wire w4;    //: /sn:0 {0}(252,278)(164,278){1}
wire w0;    //: /sn:0 {0}(318,174)(696,174)(696,241)(735,241){1}
wire w3;    //: /sn:0 {0}(251,78)(164,78){1}
wire w12;    //: /sn:0 {0}(318,126)(706,126)(706,231)(735,231){1}
wire w19;    //: /sn:0 {0}(318,442)(718,442)(718,291)(735,291){1}
wire w10;    //: /sn:0 {0}(318,279)(688,279)(688,261)(735,261){1}
wire w1;    //: /sn:0 {0}(735,221)(716,221)(716,79)(317,79){1}
wire w8;    //: /sn:0 {0}(251,173)(164,173){1}
wire w14;    //: /sn:0 {0}(318,332)(697,332)(697,271)(735,271){1}
wire w11;    //: /sn:0 {0}(252,223)(164,223){1}
wire w5;    //: /sn:0 {0}(251,125)(164,125){1}
wire w9;    //: /sn:0 {0}(251,386)(164,386){1}
//: enddecls

  //: OUT g4 (out) @(809,256) /sn:0 /tech:unit /w:[ 0 ]
  //: IN g8 (clk) @(208,512) /sn:0 /R:1 /tech:unit /w:[ 29 ]
  assign out = {w19, w6, w14, w10, w16, w0, w12, w1}; //: CONCAT g3  @(740,256) /sn:0 /w:[ 1 1 1 1 1 1 1 1 0 ] /dr:1 /tp:0 /drp:1
  FFDet g16 (.D(w4), .clk(clk), .Y(w10));   //: @(253, 269) /sz:(64, 45) /sn:0 /p:[ Li0>0 Li1>15 Ro0<0 ]
  FFDet g26 (.D(w13), .clk(clk), .Y(w19));   //: @(252, 432) /sz:(65, 45) /sn:0 /p:[ Li0>1 Li1>27 Ro0<0 ]
  FFDet g17 (.D(w9), .clk(clk), .Y(w6));   //: @(252, 377) /sz:(65, 45) /sn:0 /p:[ Li0>0 Li1>23 Ro0<0 ]
  FFDet g2 (.D(w3), .clk(clk), .Y(w1));   //: @(252, 69) /sz:(64, 45) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  //: joint g23 (clk) @(208, 410) /w:[ 22 21 -1 24 ]
  assign w3 = in[0]; //: TAP g1 @(158,78) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: joint g24 (clk) @(208, 300) /w:[ 14 13 -1 16 ]
  //: joint g18 (clk) @(208, 465) /w:[ 26 25 -1 28 ]
  //: joint g25 (clk) @(208, 355) /w:[ 18 17 -1 20 ]
  //: joint g10 (clk) @(208, 196) /w:[ 6 5 -1 8 ]
  FFDet g6 (.D(w8), .clk(clk), .Y(w0));   //: @(252, 165) /sz:(65, 43) /sn:0 /p:[ Li0>0 Li1>7 Ro0<0 ]
  FFDet g7 (.D(w11), .clk(clk), .Y(w16));   //: @(253, 214) /sz:(64, 46) /sn:0 /p:[ Li0>0 Li1>11 Ro0<0 ]
  //: joint g9 (clk) @(208, 248) /w:[ 10 9 -1 12 ]
  assign w13 = in[7]; //: TAP g22 @(158,441) /sn:0 /R:2 /w:[ 0 16 15 ] /ss:1
  assign w5 = in[1]; //: TAP g12 @(158,125) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  FFDet g5 (.D(w5), .clk(clk), .Y(w12));   //: @(252, 117) /sz:(65, 43) /sn:0 /p:[ Li0>0 Li1>3 Ro0<0 ]
  assign w11 = in[3]; //: TAP g14 @(158,223) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: joint g11 (clk) @(208, 149) /w:[ 2 1 -1 4 ]
  FFDet g19 (.D(w7), .clk(clk), .Y(w14));   //: @(253, 323) /sz:(64, 44) /sn:0 /p:[ Li0>0 Li1>19 Ro0<0 ]
  assign w9 = in[6]; //: TAP g21 @(158,386) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  assign w7 = in[5]; //: TAP g20 @(158,331) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  //: IN g0 (in) @(160,37) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  assign w4 = in[4]; //: TAP g15 @(158,278) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  assign w8 = in[2]; //: TAP g13 @(158,173) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin MUX2x4
module MUX2x4(IN1, c, IN0, OUT);
//: interface  /sz:(98, 47) /bd:[ Ti0>IN1[3:0](70/98) Ti1>IN0[3:0](30/98) Li0>c(24/47) Bo0<OUT[3:0](52/98) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output [3:0] OUT;    //: /sn:0 {0}(#:658,273)(714,273)(714,272)(736,272){1}
input [3:0] IN1;    //: /sn:0 {0}(#:91,457)(91,401){1}
//: {2}(91,400)(91,293){3}
//: {4}(91,292)(91,188){5}
//: {6}(91,187)(91,82){7}
//: {8}(91,81)(91,24)(#:-23,24){9}
input [3:0] IN0;    //: /sn:0 {0}(#:-12,0)(166,0)(166,50){1}
//: {2}(166,51)(166,161){3}
//: {4}(166,162)(166,261){5}
//: {6}(166,262)(166,368){7}
//: {8}(166,369)(166,458){9}
input c;    //: /sn:0 {0}(71,470)(291,470)(291,438){1}
//: {2}(293,436)(412,436)(412,416){3}
//: {4}(291,434)(291,336){5}
//: {6}(293,334)(412,334)(412,308){7}
//: {8}(291,332)(291,222){9}
//: {10}(293,220)(411,220)(411,206){11}
//: {12}(291,218)(291,111)(410,111)(410,98){13}
wire w13;    //: /sn:0 {0}(360,290)(103,290)(103,293)(95,293){1}
wire w7;    //: /sn:0 {0}(457,172)(590,172)(590,268)(652,268){1}
wire w4;    //: /sn:0 {0}(361,157)(178,157)(178,162)(170,162){1}
wire w3;    //: /sn:0 {0}(456,64)(641,64)(641,258)(652,258){1}
wire w0;    //: /sn:0 {0}(362,80)(103,80)(103,82)(95,82){1}
wire w12;    //: /sn:0 {0}(360,259)(178,259)(178,262)(170,262){1}
wire w1;    //: /sn:0 {0}(362,49)(178,49)(178,51)(170,51){1}
wire w8;    //: /sn:0 {0}(359,367)(178,367)(178,369)(170,369){1}
wire w11;    //: /sn:0 {0}(652,288)(536,288)(536,382)(460,382){1}
wire w15;    //: /sn:0 {0}(459,274)(475,274)(475,278)(652,278){1}
wire w5;    //: /sn:0 {0}(361,188)(95,188){1}
wire w9;    //: /sn:0 {0}(359,398)(103,398)(103,401)(95,401){1}
//: enddecls

  myMUX2 g4 (.a(w12), .b(w13), .c(c), .out(w15));   //: @(361, 245) /sz:(97, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>7 Ro0<0 ]
  myMUX2 g3 (.a(w8), .b(w9), .c(c), .out(w11));   //: @(360, 353) /sz:(99, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>3 Ro0<1 ]
  //: IN g17 (IN1) @(-25,24) /sn:0 /w:[ 9 ]
  //: IN g26 (c) @(69,470) /sn:0 /w:[ 0 ]
  myMUX2 g2 (.a(w4), .b(w5), .c(c), .out(w7));   //: @(362, 143) /sz:(94, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>11 Ro0<0 ]
  //: IN g1 (IN0) @(-14,0) /sn:0 /w:[ 0 ]
  assign w0 = IN1[0]; //: TAP g18 @(89,82) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1
  assign w4 = IN0[1]; //: TAP g10 @(164,162) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  assign w1 = IN0[0]; //: TAP g9 @(164,51) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: OUT g35 (OUT) @(733,272) /sn:0 /w:[ 1 ]
  //: joint g31 (c) @(291, 436) /w:[ 2 4 -1 1 ]
  //: joint g33 (c) @(291, 220) /w:[ 10 12 -1 9 ]
  assign w8 = IN0[3]; //: TAP g12 @(164,369) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  assign OUT = {w11, w15, w7, w3}; //: CONCAT g34  @(657,273) /sn:0 /w:[ 0 0 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign w12 = IN0[2]; //: TAP g11 @(164,262) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  assign w5 = IN1[1]; //: TAP g19 @(89,188) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  assign w9 = IN1[3]; //: TAP g21 @(89,401) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:1
  assign w13 = IN1[2]; //: TAP g20 @(89,293) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  //: joint g32 (c) @(291, 334) /w:[ 6 8 -1 5 ]
  myMUX2 g0 (.a(w1), .b(w0), .c(c), .out(w3));   //: @(363, 35) /sz:(92, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>13 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUX2x8
module MUX2x8(IN1, c, IN0, OUT);
//: interface  /sz:(47, 111) /bd:[ Li0>IN1[7:0](25/111) Li1>IN0[7:0](82/111) Bi0>c(11/47) Ro0<OUT[7:0](53/111) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output [7:0] OUT;    //: /sn:0 {0}(#:816,422)(940,422)(940,408)(955,408){1}
input [7:0] IN1;    //: /sn:0 {0}(#:241,929)(241,887){1}
//: {2}(241,886)(241,799){3}
//: {4}(241,798)(241,713){5}
//: {6}(241,712)(241,625){7}
//: {8}(241,624)(241,535){9}
//: {10}(241,534)(241,477)(242,477)(242,439){11}
//: {12}(242,438)(242,356){13}
//: {14}(242,355)(242,268){15}
//: {16}(242,267)(242,223)(#:131,223){17}
input [7:0] IN0;    //: /sn:0 {0}(#:162,200)(317,200)(317,229){1}
//: {2}(317,230)(317,324){3}
//: {4}(317,325)(317,407){5}
//: {6}(317,408)(317,503){7}
//: {8}(317,504)(317,593){9}
//: {10}(317,594)(317,634)(318,634)(318,681){11}
//: {12}(318,682)(318,767){13}
//: {14}(318,768)(318,795)(317,795)(317,858){15}
//: {16}(317,859)(317,949){17}
input c;    //: /sn:0 {0}(556,374)(556,388)(445,388){1}
//: {2}(443,386)(443,303)(556,303)(556,290){3}
//: {4}(443,390)(443,445)(442,445)(442,481){5}
//: {6}(444,483)(557,483)(557,457){7}
//: {8}(442,485)(442,522)(441,522)(441,571){9}
//: {10}(443,573)(557,573)(557,553){11}
//: {12}(441,575)(441,652){13}
//: {14}(443,654)(556,654)(556,643){15}
//: {16}(441,656)(441,740){17}
//: {18}(443,742)(555,742)(555,731){19}
//: {20}(441,744)(441,832){21}
//: {22}(443,834)(553,834)(553,817){23}
//: {24}(441,836)(441,909){25}
//: {26}(443,911)(554,911)(554,905){27}
//: {28}(441,913)(441,956)(207,956){29}
wire w13;    //: /sn:0 {0}(511,439)(246,439){1}
wire w16;    //: /sn:0 {0}(505,768)(322,768){1}
wire w7;    //: /sn:0 {0}(607,340)(776,340)(776,397)(810,397){1}
wire w4;    //: /sn:0 {0}(511,325)(321,325){1}
wire w25;    //: /sn:0 {0}(505,713)(245,713){1}
wire w0;    //: /sn:0 {0}(511,268)(246,268){1}
wire w3;    //: /sn:0 {0}(607,248)(799,248)(799,387)(810,387){1}
wire w29;    //: /sn:0 {0}(507,625)(245,625){1}
wire w12;    //: /sn:0 {0}(511,408)(321,408){1}
wire w19;    //: /sn:0 {0}(608,783)(749,783)(749,447)(810,447){1}
wire w23;    //: /sn:0 {0}(609,872)(768,872)(768,457)(810,457){1}
wire w21;    //: /sn:0 {0}(506,887)(245,887){1}
wire w24;    //: /sn:0 {0}(505,682)(322,682){1}
wire w1;    //: /sn:0 {0}(511,230)(321,230){1}
wire w31;    //: /sn:0 {0}(810,427)(727,427)(727,526)(714,526)(714,609)(612,609){1}
wire w32;    //: /sn:0 {0}(506,858)(330,858)(330,859)(321,859){1}
wire w8;    //: /sn:0 {0}(509,504)(321,504){1}
wire w17;    //: /sn:0 {0}(505,799)(245,799){1}
wire w27;    //: /sn:0 {0}(810,437)(732,437)(732,697)(611,697){1}
wire w28;    //: /sn:0 {0}(507,594)(321,594){1}
wire w11;    //: /sn:0 {0}(810,417)(719,417)(719,519)(610,519){1}
wire w15;    //: /sn:0 {0}(608,423)(713,423)(713,407)(810,407){1}
wire w5;    //: /sn:0 {0}(511,356)(246,356){1}
wire w9;    //: /sn:0 {0}(509,535)(245,535){1}
//: enddecls

  myMUX2 g4 (.a(w12), .b(w13), .c(c), .out(w15));   //: @(512, 394) /sz:(95, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>7 Ro0<0 ]
  myMUX2 g8 (.a(w28), .b(w29), .c(c), .out(w31));   //: @(508, 580) /sz:(103, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>15 Ro0<1 ]
  myMUX2 g3 (.a(w8), .b(w9), .c(c), .out(w11));   //: @(510, 490) /sz:(99, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>11 Ro0<1 ]
  assign w32 = IN0[7]; //: TAP g16 @(315,859) /sn:0 /R:2 /w:[ 1 16 15 ] /ss:1
  //: IN g17 (IN1) @(129,223) /sn:0 /w:[ 17 ]
  //: IN g26 (c) @(205,956) /sn:0 /w:[ 29 ]
  myMUX2 g2 (.a(w4), .b(w5), .c(c), .out(w7));   //: @(512, 311) /sz:(94, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>0 Ro0<0 ]
  assign w25 = IN1[5]; //: TAP g23 @(239,713) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  //: joint g30 (c) @(441, 654) /w:[ 14 13 -1 16 ]
  //: IN g1 (IN0) @(160,200) /sn:0 /w:[ 0 ]
  assign w17 = IN1[6]; //: TAP g24 @(239,799) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  //: joint g29 (c) @(441, 742) /w:[ 18 17 -1 20 ]
  assign w0 = IN1[0]; //: TAP g18 @(240,268) /sn:0 /R:2 /w:[ 1 15 16 ] /ss:1
  assign w4 = IN0[1]; //: TAP g10 @(315,325) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  assign w21 = IN1[7]; //: TAP g25 @(239,887) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:1
  myMUX2 g6 (.a(w32), .b(w21), .c(c), .out(w23));   //: @(507, 845) /sz:(101, 59) /sn:0 /p:[ Li0>0 Li1>0 Bi0>27 Ro0<0 ]
  myMUX2 g7 (.a(w24), .b(w25), .c(c), .out(w27));   //: @(506, 668) /sz:(104, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>19 Ro0<1 ]
  assign w1 = IN0[0]; //: TAP g9 @(315,230) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: OUT g35 (OUT) @(952,408) /sn:0 /w:[ 1 ]
  assign w29 = IN1[4]; //: TAP g22 @(239,625) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1
  //: joint g31 (c) @(441, 573) /w:[ 10 9 -1 12 ]
  //: joint g33 (c) @(443, 388) /w:[ 1 2 -1 4 ]
  assign w8 = IN0[3]; //: TAP g12 @(315,504) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: joint g28 (c) @(441, 834) /w:[ 22 21 -1 24 ]
  assign OUT = {w23, w19, w27, w31, w11, w15, w7, w3}; //: CONCAT g34  @(815,422) /sn:0 /w:[ 0 1 1 0 0 0 1 1 1 ] /dr:1 /tp:0 /drp:1
  myMUX2 g5 (.a(w16), .b(w17), .c(c), .out(w19));   //: @(506, 754) /sz:(101, 62) /sn:0 /p:[ Li0>0 Li1>0 Bi0>23 Ro0<0 ]
  assign w12 = IN0[2]; //: TAP g11 @(315,408) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  assign w24 = IN0[5]; //: TAP g14 @(316,682) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  assign w5 = IN1[1]; //: TAP g19 @(240,356) /sn:0 /R:2 /w:[ 1 13 14 ] /ss:1
  assign w9 = IN1[3]; //: TAP g21 @(239,535) /sn:0 /R:2 /w:[ 1 9 10 ] /ss:1
  assign w13 = IN1[2]; //: TAP g20 @(240,439) /sn:0 /R:2 /w:[ 1 11 12 ] /ss:1
  //: joint g32 (c) @(442, 483) /w:[ 6 5 -1 8 ]
  myMUX2 g0 (.a(w1), .b(w0), .c(c), .out(w3));   //: @(512, 213) /sz:(94, 76) /sn:0 /p:[ Li0>0 Li1>0 Bi0>3 Ro0<0 ]
  assign w16 = IN0[6]; //: TAP g15 @(316,768) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  //: joint g27 (c) @(441, 911) /w:[ 26 25 -1 28 ]
  assign w28 = IN0[4]; //: TAP g13 @(315,594) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin MUL_ADD
module MUL_ADD(clk, D, C, B, c, S, A);
//: interface  /sz:(98, 49) /bd:[ Ti0>A[3:0](18/98) Ti1>B[3:0](39/98) Ti2>C[3:0](60/98) Ti3>D[3:0](78/98) Li0>c(16/49) Li1>clk(33/49) Bo0<S[7:0](48/98) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] B;    //: /sn:0 {0}(#:686,74)(686,99){1}
input [3:0] A;    //: /sn:0 {0}(#:644,74)(644,99){1}
input clk;    //: /sn:0 {0}(695,368)(695,328)(479,328){1}
supply0 w14;    //: /sn:0 {0}(792,293)(808,293){1}
input [3:0] C;    //: /sn:0 {0}(#:743,78)(743,99){1}
input [3:0] D;    //: /sn:0 {0}(#:785,79)(785,99){1}
output [7:0] S;    //: /sn:0 {0}(#:723,197)(723,187)(#:585,187)(585,440)(724,440){1}
//: {2}(726,438)(726,418){3}
//: {4}(726,442)(#:726,510){5}
input c;    //: /sn:0 {0}(636,209)(484,209){1}
wire [7:0] MUL2;    //: /sn:0 {0}(#:763,271)(763,141){1}
wire [7:0] SOMMAinterno;    //: /sn:0 {0}(726,368)(#:726,317){1}
wire [7:0] MUX;    //: /sn:0 {0}(#:695,271)(#:695,246){1}
wire [7:0] MUL1;    //: /sn:0 {0}(#:666,141)(#:666,197){1}
wire w79;    //: /sn:0 {0}(665,295)(650,295){1}
//: enddecls

  //: IN g4 (clk) @(477,328) /sn:0 /tech:unit /w:[ 1 ]
  //: IN g3 (D) @(785,77) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  //: IN g2 (C) @(743,76) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  //: IN g1 (B) @(686,72) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  //: joint g6 (S) @(726, 440) /w:[ -1 2 1 4 ]
  //: IN g7 (c) @(482,209) /sn:0 /tech:unit /w:[ 1 ]
  //: GROUND g59 (w14) @(814,293) /sn:0 /R:1 /w:[ 1 ]
  MUX2x8 g36 (.IN0(MUL1), .IN1(S), .c(c), .OUT(MUX));   //: @(638, 198) /sz:(111, 47) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Bo0<1 ]
  MUL4 g14 (.A(A), .B(B), .S(MUL1));   //: @(617, 100) /sz:(92, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 ]
  //: OUT g5 (S) @(726,507) /sn:0 /R:3 /tech:unit /w:[ 5 ]
  MUL4 g32 (.A(C), .B(D), .S(MUL2));   //: @(716, 100) /sz:(92, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]
  //: IN g0 (A) @(644,72) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  RCA8 g48 (.A(MUX), .B(MUL2), .Cin(w14), .Cout(w79), .S(SOMMAinterno));   //: @(666, 272) /sz:(125, 44) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  SReg8 g13 (.clk(clk), .in(SOMMAinterno), .out(S));   //: @(685, 369) /sz:(88, 48) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<3 ]

endmodule
//: /netlistEnd

//: /netlistBegin SReg4
module SReg4(out, clk, in);
//: interface  /sz:(106, 52) /bd:[ Ti0>clk(14/106) Ti1>in[3:0](54/106) Bo0<out[3:0](55/106) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] in;    //: /sn:0 {0}(#:12,-282)(12,-236){1}
//: {2}(12,-235)(12,-155){3}
//: {4}(12,-154)(12,-89){5}
//: {6}(12,-88)(12,-19){7}
//: {8}(12,-18)(12,48){9}
output [3:0] out;    //: /sn:0 {0}(#:408,-114)(441,-114){1}
input clk;    //: /sn:0 {0}(103,7)(59,7){1}
//: {2}(57,5)(57,-62){3}
//: {4}(59,-64)(103,-64){5}
//: {6}(57,-66)(57,-128){7}
//: {8}(59,-130)(103,-130){9}
//: {10}(57,-132)(57,-211)(103,-211){11}
//: {12}(57,9)(57,59){13}
wire w16;    //: /sn:0 {0}(169,-17)(353,-17)(353,-99)(402,-99){1}
wire w0;    //: /sn:0 {0}(170,-87)(315,-87)(315,-109)(402,-109){1}
wire w3;    //: /sn:0 {0}(103,-235)(16,-235){1}
wire w12;    //: /sn:0 {0}(170,-153)(314,-153)(314,-119)(402,-119){1}
wire w1;    //: /sn:0 {0}(402,-129)(350,-129)(350,-234)(169,-234){1}
wire w8;    //: /sn:0 {0}(103,-88)(16,-88){1}
wire w11;    //: /sn:0 {0}(103,-18)(16,-18){1}
wire w5;    //: /sn:0 {0}(103,-154)(16,-154){1}
//: enddecls

  //: OUT g4 (out) @(438,-114) /sn:0 /tech:unit /w:[ 1 ]
  //: IN g8 (clk) @(57,61) /sn:0 /R:1 /tech:unit /w:[ 13 ]
  assign out = {w16, w0, w12, w1}; //: CONCAT g3  @(407,-114) /sn:0 /w:[ 0 1 1 1 0 ] /dr:1 /tp:1 /drp:1
  FFDet g2 (.D(w3), .clk(clk), .Y(w1));   //: @(104, -244) /sz:(64, 45) /sn:0 /p:[ Li0>0 Li1>11 Ro0<1 ]
  assign w3 = in[0]; //: TAP g1 @(10,-235) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: joint g10 (clk) @(57, -64) /w:[ 4 6 -1 3 ]
  FFDet g6 (.D(w8), .clk(clk), .Y(w0));   //: @(104, -97) /sz:(65, 45) /sn:0 /p:[ Li0>0 Li1>5 Ro0<0 ]
  FFDet g7 (.D(w11), .clk(clk), .Y(w16));   //: @(104, -27) /sz:(64, 46) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  //: joint g9 (clk) @(57, -130) /w:[ 8 10 -1 7 ]
  assign w5 = in[1]; //: TAP g12 @(10,-154) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  FFDet g5 (.D(w5), .clk(clk), .Y(w12));   //: @(104, -162) /sz:(65, 43) /sn:0 /p:[ Li0>0 Li1>9 Ro0<0 ]
  //: joint g11 (clk) @(57, 7) /w:[ 1 2 -1 12 ]
  assign w11 = in[3]; //: TAP g14 @(10,-18) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: IN g0 (in) @(12,-284) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  assign w8 = in[2]; //: TAP g13 @(10,-88) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin FA
module FA(Cin, B, A, S, Cout);
//: interface  /sz:(55, 54) /bd:[ Ti0>B(39/55) Ti1>A(14/55) Ri0>Cin(25/54) Lo0<Cout(24/54) Bo0<S(26/55) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(174,202)(174,73)(254,73){1}
//: {2}(256,71)(256,50){3}
//: {4}(256,75)(256,109){5}
input A;    //: /sn:0 {0}(150,202)(150,62)(229,62){1}
//: {2}(231,60)(231,48){3}
//: {4}(231,64)(231,109){5}
input Cin;    //: /sn:0 {0}(80,202)(80,159)(165,159){1}
//: {2}(169,159)(218,159)(218,200){3}
//: {4}(167,157)(167,46){5}
output Cout;    //: /sn:0 {0}(130,310)(130,328){1}
output S;    //: /sn:0 {0}(227,248)(227,321){1}
wire w4;    //: /sn:0 {0}(139,265)(139,260)(164,260)(164,244){1}
wire w3;    //: /sn:0 {0}(116,265)(116,260)(94,260)(94,244){1}
wire w2;    //: /sn:0 {0}(105,202)(105,180)(238,180){1}
//: {2}(240,178)(240,151){3}
//: {4}(240,182)(240,200){5}
//: enddecls

  //: IN g4 (Cin) @(167,44) /sn:0 /R:3 /w:[ 5 ]
  //: joint g8 (w2) @(240, 180) /w:[ -1 2 1 4 ]
  //: IN g3 (B) @(256,48) /sn:0 /R:3 /w:[ 3 ]
  //: IN g2 (A) @(231,46) /sn:0 /R:3 /w:[ 3 ]
  myEXOR g1 (.B(Cin), .A(w2), .out(S));   //: @(200, 201) /sz:(54, 46) /R:3 /sn:0 /p:[ Ti0>3 Ti1>5 Bo0<0 ]
  myNAND g10 (.in2(A), .in1(B), .out(w4));   //: @(134, 203) /sz:(56, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  //: OUT g6 (S) @(227,318) /sn:0 /R:3 /w:[ 1 ]
  myNAND g7 (.in2(Cin), .in1(w2), .out(w3));   //: @(63, 203) /sz:(58, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  //: joint g9 (Cin) @(167, 159) /w:[ 2 4 1 -1 ]
  //: joint g12 (B) @(256, 73) /w:[ -1 2 1 4 ]
  //: OUT g5 (Cout) @(130,325) /sn:0 /R:3 /w:[ 1 ]
  //: joint g11 (A) @(231, 62) /w:[ -1 2 1 4 ]
  myEXOR g0 (.B(A), .A(B), .out(w2));   //: @(213, 110) /sz:(54, 40) /R:2 /sn:0 /p:[ Ti0>5 Ti1>5 Bo0<3 ]
  myNAND g13 (.in2(w3), .in1(w4), .out(Cout));   //: @(101, 266) /sz:(53, 43) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUL_SUB
module MUL_SUB(Cout, S, A, C, B);
//: interface  /sz:(164, 68) /bd:[ Ti0>A[7:0](80/164) Ri0>B[3:0](16/68) Ri1>C[3:0](53/68) Lo0<Cout(35/68) Bo0<S[7:0](81/164) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
supply1 w7;    //: /sn:0 {0}(589,490)(598,490)(598,454){1}
input [3:0] B;    //: /sn:0 {0}(#:521,311)(#:521,355){1}
input [7:0] A;    //: /sn:0 {0}(513,467)(513,441)(436,441)(#:436,313){1}
output Cout;    //: /sn:0 {0}(491,490)(379,490){1}
input [3:0] C;    //: /sn:0 {0}(#:563,310)(#:563,355){1}
output [7:0] S;    //: /sn:0 {0}(#:535,509)(535,545)(383,545){1}
wire [7:0] w19;    //: /sn:0 {0}(#:543,397)(543,467){1}
//: enddecls

  //: OUT g4 (Cout) @(382,490) /sn:0 /R:2 /tech:unit /w:[ 1 ]
  //: VDD g16 (w7) @(609,454) /sn:0 /tech:unit /w:[ 1 ]
  //: OUT g3 (S) @(386,545) /sn:0 /R:2 /tech:unit /w:[ 1 ]
  //: IN g2 (A) @(436,311) /sn:0 /R:3 /tech:unit /w:[ 1 ]
  MUL4 g91 (.A(B), .B(C), .S(w19));   //: @(494, 356) /sz:(92, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 ]
  //: IN g1 (C) @(563,308) /sn:0 /R:3 /tech:unit /w:[ 0 ]
  SUB8 g15 (.A(A), .B(w19), .Cin(w7), .Cout(Cout), .S(S));   //: @(492, 468) /sz:(96, 40) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: IN g0 (B) @(521,309) /sn:0 /R:3 /tech:unit /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUL4
module MUL4(B, S, A);
//: interface  /sz:(92, 40) /bd:[ Ti0>B[3:0](69/92) Ti1>A[3:0](27/92) Bo0<S[7:0](49/92) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] B;    //: /sn:0 {0}(#:721,-464)(676,-464){1}
//: {2}(675,-464)(411,-464){3}
//: {4}(410,-464)(148,-464){5}
//: {6}(147,-464)(-68,-464){7}
//: {8}(-69,-464)(-216,-464){9}
input [3:0] A;    //: /sn:0 {0}(#:445,-514)(449,-514){1}
//: {2}(450,-514)(519,-514){3}
//: {4}(520,-514)(586,-514){5}
//: {6}(587,-514)(656,-514){7}
//: {8}(657,-514)(#:723,-514){9}
output [7:0] S;    //: /sn:0 {0}(#:71,167)(71,204){1}
wire w13;    //: /sn:0 {0}(-140,-394)(-140,-435)(72,-435){1}
//: {2}(76,-435)(320,-435){3}
//: {4}(324,-435)(585,-435){5}
//: {6}(587,-437)(587,-510){7}
//: {8}(587,-433)(587,-397){9}
//: {10}(322,-433)(322,-394){11}
//: {12}(74,-433)(74,-394){13}
wire w16;    //: /sn:0 {0}(-87,-394)(-87,-417)(127,-417){1}
//: {2}(131,-417)(389,-417){3}
//: {4}(393,-417)(655,-417){5}
//: {6}(657,-419)(657,-510){7}
//: {8}(657,-415)(657,-399){9}
//: {10}(391,-415)(391,-396){11}
//: {12}(129,-415)(129,-394){13}
wire w7;    //: /sn:0 {0}(-245,-394)(-245,-451)(-32,-451){1}
//: {2}(-28,-451)(183,-451){3}
//: {4}(187,-451)(448,-451){5}
//: {6}(450,-453)(450,-510){7}
//: {8}(450,-449)(450,-397){9}
//: {10}(185,-449)(185,-394){11}
//: {12}(-30,-449)(-30,-394){13}
wire w34;    //: /sn:0 {0}(218,11)(178,11)(178,-23)(146,-23)(146,-13){1}
wire w25;    //: /sn:0 {0}(166,-214)(218,-214){1}
wire w4;    //: /sn:0 {0}(-17,-352)(-17,-281)(24,-281)(24,-241){1}
wire w109;    //: /sn:0 {0}(36,161)(36,123)(-146,123)(-146,13)(-123,13){1}
wire w22;    //: /sn:0 {0}(32,-353)(32,-292)(112,-292)(112,-240){1}
wire w36;    //: /sn:0 {0}(76,161)(76,113)(254,113)(254,41){1}
wire w0;    //: /sn:0 {0}(-194,-394)(-194,-442)(21,-442){1}
//: {2}(25,-442)(253,-442){3}
//: {4}(257,-442)(518,-442){5}
//: {6}(520,-444)(520,-510){7}
//: {8}(520,-440)(520,-399){9}
//: {10}(255,-440)(255,-396){11}
//: {12}(23,-440)(23,-395){13}
wire w20;    //: /sn:0 {0}(264,-354)(264,-327)(236,-327)(236,-239){1}
wire w60;    //: /sn:0 {0}(86,161)(86,126)(379,126)(379,-63){1}
wire w29;    //: /sn:0 {0}(-78,-352)(-78,-32)(234,-32)(234,-17){1}
wire w37;    //: /sn:0 {0}(479,-212)(417,-212){1}
wire w12;    //: /sn:0 {0}(46,-215)(94,-215){1}
wire w19;    //: /sn:0 {0}(7,-183)(7,-59)(-4,-59)(-4,-11){1}
wire w18;    //: /sn:0 {0}(204,-394)(204,-424)(272,-424){1}
//: {2}(276,-424)(339,-424){3}
//: {4}(343,-424)(409,-424){5}
//: {6}(411,-426)(411,-460){7}
//: {8}(411,-422)(411,-409)(410,-409)(410,-396){9}
//: {10}(341,-422)(341,-394){11}
//: {12}(274,-422)(274,-396){13}
wire w23;    //: /sn:0 {0}(194,-352)(194,-291)(144,-291)(144,-240){1}
wire w10;    //: /sn:0 {0}(-185,-352)(-185,-271)(-9,-271)(-9,-241){1}
wire w70;    //: /sn:0 {0}(268,-17)(268,-47)(253,-47)(253,-63){1}
wire w54;    //: /sn:0 {0}(343,-93)(290,-93){1}
wire w24;    //: /sn:0 {0}(-11,-394)(-11,-426)(40,-426){1}
//: {2}(44,-426)(91,-426){3}
//: {4}(95,-426)(146,-426){5}
//: {6}(148,-428)(148,-460){7}
//: {8}(148,-424)(148,-394){9}
//: {10}(93,-424)(93,-394){11}
//: {12}(42,-424)(42,-395){13}
wire w31;    //: /sn:0 {0}(131,-184)(131,-156)(147,-156)(147,-120){1}
wire w1;    //: /sn:0 {0}(469,-397)(469,-431)(537,-431){1}
//: {2}(541,-431)(604,-431){3}
//: {4}(608,-431)(674,-431){5}
//: {6}(676,-433)(676,-460){7}
//: {8}(676,-429)(676,-399){9}
//: {10}(606,-429)(606,-397){11}
//: {12}(539,-429)(539,-399){13}
wire w104;    //: /sn:0 {0}(-51,14)(-23,14){1}
wire w32;    //: /sn:0 {0}(359,-122)(359,-155)(318,-155)(318,-278)(138,-278)(138,-352){1}
wire w8;    //: /sn:0 {0}(459,-355)(459,-316)(267,-316)(267,-239){1}
wire w110;    //: /sn:0 {0}(46,161)(46,104)(-89,104)(-89,44){1}
wire w46;    //: /sn:0 {0}(29,-11)(29,-95)(96,-95){1}
wire w89;    //: /sn:0 {0}(251,-183)(251,-155)(268,-155)(268,-119){1}
wire w27;    //: /sn:0 {0}(-226,-394)(-226,-422)(-177,-422){1}
//: {2}(-173,-422)(-123,-422){3}
//: {4}(-119,-422)(-70,-422){5}
//: {6}(-68,-424)(-68,-460){7}
//: {8}(-68,-420)(-68,-394){9}
//: {10}(-121,-420)(-121,-394){11}
//: {12}(-175,-420)(-175,-394){13}
wire w17;    //: /sn:0 {0}(400,-354)(400,-297)(488,-297)(488,-254)(494,-254)(494,-242){1}
wire w35;    //: /sn:0 {0}(-236,-352)(-236,-27)(-105,-27)(-105,-12){1}
wire w28;    //: /sn:0 {0}(331,-352)(331,-267)(362,-267)(362,-239){1}
wire w45;    //: /sn:0 {0}(169,-94)(219,-94){1}
wire w2;    //: /sn:0 {0}(666,-357)(666,142)(106,142)(106,161){1}
wire w41;    //: /sn:0 {0}(-131,-352)(-131,-134)(115,-134)(115,-120){1}
wire w11;    //: /sn:0 {0}(529,-357)(529,-267)(395,-267)(395,-239){1}
wire w47;    //: /sn:0 {0}(132,-64)(132,-22)(112,-22)(112,-13){1}
wire w105;    //: /sn:0 {0}(56,161)(56,81)(12,81)(12,47){1}
wire w15;    //: /sn:0 {0}(-73,-12)(-73,-25)(-94,-25)(-94,-216)(-28,-216){1}
wire w38;    //: /sn:0 {0}(83,-352)(83,-307)(200,-307)(200,-177)(237,-177)(237,-119){1}
wire w92;    //: /sn:0 {0}(517,-180)(517,132)(96,132)(96,161){1}
wire w5;    //: /sn:0 {0}(596,-355)(596,-296)(536,-296)(536,-254)(528,-254)(528,-242){1}
wire w43;    //: /sn:0 {0}(393,-122)(393,-140)(380,-140)(380,-179){1}
wire w100;    //: /sn:0 {0}(66,161)(66,104)(132,104)(132,44){1}
wire w99;    //: /sn:0 {0}(52,15)(96,15){1}
wire w40;    //: /sn:0 {0}(288,-213)(343,-213){1}
//: enddecls

  FA g116 (.A(w28), .B(w11), .Cin(w37), .Cout(w40), .S(w43));   //: @(344, -238) /sz:(72, 58) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  myAND g4 (.in1(w1), .in2(w13), .out(w5));   //: @(575, -396) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>11 Ti1>9 Bo0<0 ]
  myAND g8 (.in1(w18), .in2(w16), .out(w17));   //: @(379, -395) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>9 Ti1>11 Bo0<0 ]
  myAND g16 (.in1(w27), .in2(w13), .out(w41));   //: @(-152, -393) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>11 Ti1>0 Bo0<0 ]
  assign w16 = A[0]; //: TAP g3 @(657,-516) /sn:0 /R:1 /w:[ 7 7 8 ] /ss:1
  //: joint g109 (w0) @(23, -442) /w:[ 2 -1 1 12 ]
  myAND g17 (.in1(w27), .in2(w0), .out(w10));   //: @(-206, -393) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>13 Ti1>0 Bo0<0 ]
  assign w18 = B[1]; //: TAP g26 @(411,-466) /sn:0 /R:1 /w:[ 7 4 3 ] /ss:1
  myAND g2 (.in1(w1), .in2(w16), .out(w2));   //: @(645, -398) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>9 Ti1>9 Bo0<0 ]
  //: joint g23 (w1) @(676, -431) /w:[ -1 6 5 8 ]
  //: joint g30 (w27) @(-121, -422) /w:[ 4 -1 3 10 ]
  //: joint g104 (w13) @(587, -435) /w:[ -1 6 5 8 ]
  //: IN g1 (B) @(723,-464) /sn:0 /R:2 /tech:unit /w:[ 0 ]
  //: joint g24 (w1) @(606, -431) /w:[ 4 -1 3 10 ]
  //: joint g111 (w7) @(185, -451) /w:[ 4 -1 3 10 ]
  //: joint g110 (w7) @(450, -451) /w:[ -1 6 5 8 ]
  //: joint g29 (w27) @(-68, -422) /w:[ -1 6 5 8 ]
  myAND g18 (.in1(w24), .in2(w7), .out(w4));   //: @(-42, -393) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>13 Bo0<0 ]
  FA g70 (.B(w46), .A(w19), .Cin(w99), .Cout(w104), .S(w105));   //: @(-22, -10) /sz:(73, 56) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  //: joint g103 (w18) @(274, -424) /w:[ 2 -1 1 12 ]
  myAND g10 (.in1(w18), .in2(w7), .out(w23));   //: @(173, -393) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>11 Bo0<0 ]
  //: joint g25 (w1) @(539, -431) /w:[ 2 -1 1 12 ]
  //: joint g107 (w0) @(520, -442) /w:[ -1 6 5 8 ]
  assign S = {w109, w110, w105, w100, w36, w60, w92, w2}; //: CONCAT g72  @(71,166) /sn:0 /R:3 /tech:unit /w:[ 0 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  myAND g6 (.in1(w1), .in2(w0), .out(w11));   //: @(508, -398) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>13 Ti1>9 Bo0<0 ]
  FA g35 (.A(w41), .B(w31), .Cin(w45), .Cout(w46), .S(w47));   //: @(97, -119) /sz:(71, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  myAND g7 (.in1(w18), .in2(w13), .out(w28));   //: @(310, -393) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>11 Ti1>11 Bo0<0 ]
  myAND g9 (.in1(w18), .in2(w0), .out(w20));   //: @(243, -395) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>13 Ti1>11 Bo0<0 ]
  //: OUT g73 (S) @(71,201) /sn:0 /R:3 /tech:unit /w:[ 1 ]
  //: joint g102 (w18) @(341, -424) /w:[ 4 -1 3 10 ]
  assign w7 = A[3]; //: TAP g22 @(450,-516) /sn:0 /R:1 /w:[ 7 1 2 ] /ss:1
  //: joint g31 (w27) @(-175, -422) /w:[ 2 -1 1 12 ]
  FA g71 (.B(w15), .A(w35), .Cin(w104), .Cout(w109), .S(w110));   //: @(-122, -11) /sz:(70, 54) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  //: joint g99 (w16) @(391, -417) /w:[ 4 -1 3 10 ]
  FA g36 (.A(w38), .B(w89), .Cin(w54), .Cout(w45), .S(w70));   //: @(220, -118) /sz:(69, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  //: joint g33 (w24) @(93, -426) /w:[ 4 -1 3 10 ]
  //: joint g108 (w0) @(255, -442) /w:[ 4 -1 3 10 ]
  myAND g12 (.in1(w27), .in2(w16), .out(w29));   //: @(-99, -393) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>9 Ti1>0 Bo0<0 ]
  //: joint g106 (w13) @(74, -435) /w:[ 2 -1 1 12 ]
  assign w27 = B[3]; //: TAP g28 @(-68,-466) /sn:0 /R:1 /w:[ 7 8 7 ] /ss:1
  //: joint g34 (w24) @(42, -426) /w:[ 2 -1 1 12 ]
  HA g46 (.B(w34), .A(w47), .Cout(w99), .S(w100));   //: @(97, -12) /sz:(72, 55) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  myAND g5 (.in1(w1), .in2(w7), .out(w8));   //: @(438, -396) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>9 Bo0<0 ]
  myAND g11 (.in1(w24), .in2(w0), .out(w22));   //: @(11, -394) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>13 Ti1>13 Bo0<0 ]
  myAND g14 (.in1(w27), .in2(w7), .out(w35));   //: @(-257, -393) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  //: joint g112 (w7) @(-30, -451) /w:[ 2 -1 1 12 ]
  FA g117 (.A(w20), .B(w8), .Cin(w40), .Cout(w25), .S(w89));   //: @(219, -238) /sz:(68, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g114 (.A(w22), .B(w23), .Cin(w25), .Cout(w12), .S(w31));   //: @(95, -239) /sz:(70, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w1 = B[0]; //: TAP g19 @(676,-466) /sn:0 /R:1 /w:[ 7 2 1 ] /ss:1
  assign w0 = A[2]; //: TAP g21 @(520,-516) /sn:0 /R:1 /w:[ 7 3 4 ] /ss:1
  HA g115 (.A(w17), .B(w5), .Cout(w37), .S(w92));   //: @(480, -241) /sz:(71, 60) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  assign w13 = A[1]; //: TAP g20 @(587,-516) /sn:0 /R:1 /w:[ 7 5 6 ] /ss:1
  //: joint g32 (w24) @(148, -426) /w:[ -1 6 5 8 ]
  FA g113 (.A(w10), .B(w4), .Cin(w12), .Cout(w15), .S(w19));   //: @(-27, -240) /sz:(72, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g105 (w13) @(322, -435) /w:[ 4 -1 3 10 ]
  //: joint g100 (w16) @(129, -417) /w:[ 2 -1 1 12 ]
  //: joint g97 (w16) @(657, -417) /w:[ -1 6 5 8 ]
  HA g38 (.A(w29), .B(w70), .Cout(w34), .S(w36));   //: @(219, -16) /sz:(73, 56) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<1 ]
  //: joint g101 (w18) @(411, -424) /w:[ -1 6 5 8 ]
  //: IN g0 (A) @(725,-514) /sn:0 /R:2 /tech:unit /w:[ 9 ]
  myAND g15 (.in1(w24), .in2(w13), .out(w38));   //: @(62, -393) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>11 Ti1>13 Bo0<0 ]
  assign w24 = B[2]; //: TAP g27 @(148,-466) /sn:0 /R:1 /w:[ 7 6 5 ] /ss:1
  HA g37 (.A(w32), .B(w43), .Cout(w54), .S(w60));   //: @(344, -121) /sz:(72, 57) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<1 ]
  myAND g13 (.in1(w24), .in2(w16), .out(w32));   //: @(117, -393) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>9 Ti1>13 Bo0<1 ]

endmodule
//: /netlistEnd

